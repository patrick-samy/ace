module control_store(input[2:0]  address,
                     output[4:0] instruction);

    mux

endmodule
