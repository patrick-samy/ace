module micro_dispatcher(input[3:0]  opcode,
                        output[2:0] start_address);

endmodule
